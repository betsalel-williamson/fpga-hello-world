module hello_world ();

  initial begin
    $display("Hello, SystemVerilog!");
    $finish;
  end

endmodule
